library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity EntityName_TB is
end entity;

architecture test of EntityName_TB is
	
	component EntityName
		generic(
				word_size: integer;
				entries: integer);	
		port(   
				clk: in std_logic;
				rst: in std_logic;
				en: in std_logic;
				go: in std_logic;
				done: out std_logic;
				readnotwrite: in std_logic; 
				address: in std_logic_vector(word_size - 1 downto 0);
				data_in: in std_logic_vector(word_size - 1 downto 0);  
				data_out: out std_logic_vector(word_size - 1 downto 0));
	end component;

	signal clk_i : std_logic := '1';
	signal rst_i : std_logic;
	signal en_i : std_logic := '0';
	signal go_i : std_logic := '0';
	signal done_i : std_logic := '0';
	signal readnotwrite_i : std_logic := '0';
	signal address_i : std_logic_vector(8 - 1 downto 0);
	signal data_in_i : std_logic_vector(8 - 1 downto 0);
	signal data_out_i : std_logic_vector(8 - 1 downto 0);

	type resultArray is array (0 to 512 - 1) of integer;
	constant result_address_vector : resultArray := (256, 257, 258, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 286, 287, 288, 289, 290, 291, 292, 293, 294, 295, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 316, 317, 318, 319, 320, 321, 322, 323, 324, 325, 326, 327, 328, 329, 330, 331, 332, 333, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 352, 353, 354, 355, 356, 357, 358, 359, 360, 361, 362, 363, 364, 365, 366, 367, 368, 369, 370, 371, 372, 373, 374, 375, 376, 377, 378, 379, 380, 381, 382, 383, 384, 385, 386, 387, 388, 389, 390, 391, 392, 393, 394, 395, 396, 397, 398, 399, 400, 401, 402, 403, 404, 405, 406, 407, 408, 409, 410, 411, 412, 413, 414, 415, 416, 417, 418, 419, 420, 421, 422, 423, 424, 425, 426, 427, 428, 429, 430, 431, 432, 433, 434, 435, 436, 437, 438, 439, 440, 441, 442, 443, 444, 445, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 460, 461, 462, 463, 464, 465, 466, 467, 468, 469, 470, 471, 472, 473, 474, 475, 476, 477, 478, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 496, 497, 498, 499, 500, 501, 502, 503, 504, 505, 506, 507, 508, 509, 510, 511, 512, 514, 518, 523, 530, 538, 548, 559, 572, 586, 602, 619, 638, 658, 680, 703, 705, 710, 718, 729, 743, 760, 780, 803, 829, 858, 890, 925, 963, 1004, 1048, 1095, 1099, 1107, 1120, 1137, 1159, 1185, 1216, 1251, 1291, 1335, 1384, 1437, 1495, 1557, 1624, 1695, 1700, 1711, 1728, 1751, 1780, 1815, 1856, 1903, 1956, 2015, 2080, 2151, 2228, 2311, 2400, 2495, 2502, 2516, 2538, 2567, 2604, 2648, 2700, 2759, 2826, 2900, 2982, 3071, 3168, 3272, 3384, 3503, 3511, 3528, 3554, 3589, 3633, 3686, 3748, 3819, 3899, 3988, 4086, 4193, 4309, 4434, 4568, 4711, 4721, 4741, 4772, 4813, 4865, 4927, 5000, 5083, 5177, 5281, 5396, 5521, 5657, 5803, 5960, 6127, 6138, 6161, 6196, 6243, 6302, 6373, 6456, 6551, 6658, 6777, 6908, 7051, 7206, 7373, 7552, 7743, 7756, 7782, 7822, 7875, 7942, 8022, 8116, 8223, 8344, 8478, 8626, 8787, 8962, 9150, 9352, 9567, 9581, 9610, 9654, 9713, 9787, 9876, 9980, 10099, 10233, 10382, 10546, 10725, 10919, 11128, 11352, 11591, 11607, 11639, 11688, 11753, 11835, 11933, 12048, 12179, 12327, 12491, 12672, 12869, 13083, 13313, 13560, 13823, 13840, 13875, 13928, 13999, 14088, 14195, 14320, 14463, 14624, 14803, 15000, 15215, 15448, 15699, 15968, 16255, 16274, 16312, 16370, 16447, 16544, 16660, 16796, 16951, 17126, 17320, 17534, 17767, 18020, 18292, 18584, 18895, 18915, 18956, 19018, 19101, 19205, 19330, 19476, 19643, 19831, 20040, 20270, 20521, 20793, 21086, 21400, 21735, 21757, 21801, 21868, 21957, 22069, 22203, 22360, 22539, 22741, 22965, 23212, 23481, 23773, 24087, 24424, 24783, 24806, 24853, 24924, 25019, 25138, 25281, 25448, 25639, 25854, 26093, 26356, 26643, 26954, 27289, 27648, 28031);
begin

	comp: EntityName generic map (word_size => 8, entries =>28032)
									port map(clk => clk_i, rst => rst_i, en => en_i, go => go_i, done => done_i, readnotwrite => readnotwrite_i, 
									address => address_i, data_in => data_in_i, data_out => data_out_i);

	clk_i <= not(clk_i) after 0.5 ns;
	
	rst_proc : process 
		begin			
			rst_i <= '1';
			wait for 512 ns;
			rst_i <= '0';
			wait;
	end process;

	cnt_proc: process(rst_i, clk_i) 
		variable cnt : integer := 0;
		variable writeOutputs : integer := 0;
		begin
			if(rst_i = '1') then
				cnt := 0;
			elsif (clk_i'event and clk_i = '1') then
				if (cnt = 28031 and done_i = '0') then
					cnt := 0;
				elsif done_i = '1' then
					cnt := 0;
					writeOutputs := 1;
				else 
					if(writeOutputs /= 1) then
						cnt := cnt + 1;
					else
						cnt := result_address_vector(cnt);
					end if;
				end if;
			end if;
			
			address_i <= std_logic_vector(to_unsigned(cnt, 8));
	end process;

	wrt_proc: process
		variable first : boolean := true;
		begin
			if first then
				wait until en_i'event and en_i = '1' and readnotwrite_i = '0';
				first := false;
			else
				wait until en_i = '1' and readnotwrite_i = '0';
			end if;
			data_in_i <= std_logic_vector(to_unsigned(0, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(2, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(3, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(4, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(5, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(6, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(7, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(8, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(9, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(10, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(11, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(12, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(13, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(14, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(15, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(16, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(17, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(18, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(19, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(20, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(21, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(22, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(23, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(24, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(25, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(26, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(27, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(28, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(29, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(30, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(31, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(32, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(33, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(34, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(35, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(36, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(37, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(38, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(39, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(40, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(41, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(42, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(43, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(44, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(45, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(46, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(47, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(48, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(49, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(50, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(51, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(52, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(53, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(54, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(55, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(56, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(57, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(58, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(59, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(60, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(61, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(62, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(63, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(64, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(65, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(66, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(67, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(68, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(69, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(70, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(71, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(72, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(73, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(74, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(75, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(76, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(77, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(78, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(79, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(80, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(81, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(82, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(83, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(84, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(85, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(86, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(87, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(88, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(89, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(90, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(91, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(92, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(93, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(94, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(95, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(96, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(97, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(98, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(99, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(100, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(101, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(102, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(103, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(104, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(105, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(106, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(107, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(108, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(109, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(110, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(111, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(112, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(113, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(114, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(115, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(116, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(117, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(118, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(119, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(120, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(121, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(122, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(123, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(124, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(125, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(126, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(127, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(128, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(129, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(130, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(131, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(132, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(133, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(134, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(135, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(136, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(137, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(138, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(139, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(140, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(141, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(142, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(143, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(144, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(145, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(146, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(147, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(148, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(149, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(150, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(151, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(152, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(153, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(154, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(155, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(156, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(157, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(158, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(159, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(160, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(161, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(162, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(163, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(164, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(165, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(166, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(167, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(168, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(169, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(170, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(171, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(172, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(173, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(174, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(175, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(176, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(177, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(178, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(179, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(180, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(181, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(182, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(183, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(184, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(185, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(186, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(187, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(188, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(189, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(190, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(191, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(192, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(193, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(194, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(195, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(196, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(197, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(198, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(199, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(200, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(201, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(202, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(203, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(204, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(205, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(206, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(207, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(208, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(209, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(210, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(211, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(212, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(213, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(214, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(215, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(216, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(217, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(218, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(219, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(220, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(221, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(222, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(223, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(224, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(225, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(226, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(227, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(228, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(229, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(230, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(231, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(232, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(233, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(234, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(235, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(236, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(237, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(238, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(239, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(240, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(241, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(242, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(243, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(244, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(245, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(246, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(247, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(248, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(249, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(250, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(251, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(252, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(253, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(254, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(255, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(256, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(257, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(258, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(259, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(260, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(261, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(262, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(263, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(264, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(265, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(266, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(267, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(268, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(269, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(270, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(271, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(272, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(273, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(274, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(275, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(276, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(277, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(278, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(279, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(280, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(281, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(282, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(283, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(284, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(285, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(286, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(287, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(288, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(289, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(290, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(291, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(292, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(293, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(294, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(295, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(296, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(297, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(298, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(299, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(300, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(301, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(302, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(303, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(304, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(305, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(306, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(307, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(308, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(309, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(310, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(311, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(312, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(313, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(314, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(315, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(316, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(317, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(318, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(319, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(320, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(321, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(322, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(323, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(324, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(325, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(326, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(327, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(328, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(329, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(330, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(331, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(332, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(333, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(334, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(335, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(336, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(337, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(338, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(339, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(340, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(341, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(342, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(343, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(344, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(345, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(346, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(347, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(348, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(349, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(350, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(351, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(352, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(353, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(354, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(355, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(356, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(357, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(358, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(359, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(360, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(361, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(362, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(363, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(364, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(365, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(366, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(367, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(368, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(369, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(370, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(371, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(372, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(373, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(374, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(375, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(376, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(377, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(378, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(379, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(380, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(381, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(382, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(383, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(384, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(385, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(386, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(387, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(388, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(389, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(390, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(391, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(392, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(393, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(394, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(395, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(396, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(397, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(398, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(399, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(400, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(401, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(402, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(403, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(404, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(405, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(406, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(407, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(408, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(409, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(410, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(411, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(412, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(413, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(414, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(415, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(416, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(417, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(418, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(419, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(420, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(421, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(422, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(423, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(424, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(425, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(426, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(427, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(428, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(429, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(430, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(431, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(432, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(433, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(434, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(435, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(436, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(437, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(438, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(439, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(440, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(441, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(442, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(443, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(444, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(445, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(446, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(447, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(448, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(449, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(450, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(451, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(452, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(453, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(454, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(455, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(456, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(457, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(458, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(459, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(460, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(461, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(462, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(463, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(464, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(465, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(466, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(467, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(468, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(469, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(470, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(471, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(472, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(473, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(474, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(475, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(476, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(477, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(478, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(479, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(480, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(481, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(482, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(483, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(484, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(485, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(486, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(487, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(488, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(489, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(490, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(491, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(492, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(493, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(494, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(495, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(496, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(497, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(498, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(499, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(500, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(501, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(502, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(503, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(504, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(505, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(506, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(507, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(508, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(509, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(510, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(511, 8));
			wait for 1 ns;		
	end process;

	en_proc: process	
		variable first : boolean := true;
		begin
			if first then
				wait for 512 ns;
				first := false;
			end if;
			en_i <= '1';
			readnotwrite_i <= '0';
			wait for 512 ns;
			en_i <= '0';
			wait until done_i'event and done_i = '0';
			en_i <= '1';
			readnotwrite_i <= '1';
			wait for 512 ns;
	end process;

	go_proc: process
		begin
			wait until en_i'event and en_i = '0';
			go_i <= '1';
			wait for 1 ns;
			go_i <= '0';	
	end process;


end test;