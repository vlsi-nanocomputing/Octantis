library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity EntityName_TB is
end entity;

architecture test of EntityName_TB is
	
	component EntityName
		generic(
				word_size: integer;
				entries: integer);	
		port(   
				clk: in std_logic;
				rst: in std_logic;
				en: in std_logic;
				go: in std_logic;
				done: out std_logic;
				readnotwrite: in std_logic; 
				address: in std_logic_vector(word_size - 1 downto 0);
				data_in: in std_logic_vector(word_size - 1 downto 0);  
				data_out: out std_logic_vector(word_size - 1 downto 0));
	end component;

	signal clk_i : std_logic := '1';
	signal rst_i : std_logic;
	signal en_i : std_logic := '0';
	signal go_i : std_logic := '0';
	signal done_i : std_logic := '0';
	signal readnotwrite_i : std_logic := '0';
	signal address_i : std_logic_vector(8 - 1 downto 0);
	signal data_in_i : std_logic_vector(8 - 1 downto 0);
	signal data_out_i : std_logic_vector(8 - 1 downto 0);

	type resultArray is array (0 to 1536 - 1) of integer;
	constant result_address_vector : resultArray := (2564, 2565, 2566, 2567, 2568, 2569, 2570, 2571, 2572, 2573, 2574, 2575, 2576, 2577, 2578, 2579, 2580, 2581, 2582, 2583, 2584, 2585, 2586, 2587, 2588, 2589, 2590, 2591, 2592, 2593, 2594, 2595, 2596, 2597, 2598, 2599, 2600, 2601, 2602, 2603, 2604, 2605, 2606, 2607, 2608, 2609, 2610, 2611, 2612, 2613, 2614, 2615, 2616, 2617, 2618, 2619, 2620, 2621, 2622, 2623, 2624, 2625, 2626, 2627, 2628, 2629, 2630, 2631, 2632, 2633, 2634, 2635, 2636, 2637, 2638, 2639, 2640, 2641, 2642, 2643, 2644, 2645, 2646, 2647, 2648, 2649, 2650, 2651, 2652, 2653, 2654, 2655, 2656, 2657, 2658, 2659, 2660, 2661, 2662, 2663, 2664, 2665, 2666, 2667, 2668, 2669, 2670, 2671, 2672, 2673, 2674, 2675, 2676, 2677, 2678, 2679, 2680, 2681, 2682, 2683, 2684, 2685, 2686, 2687, 2688, 2689, 2690, 2691, 2692, 2693, 2694, 2695, 2696, 2697, 2698, 2699, 2700, 2701, 2702, 2703, 2704, 2705, 2706, 2707, 2708, 2709, 2710, 2711, 2712, 2713, 2714, 2715, 2716, 2717, 2718, 2719, 2720, 2721, 2722, 2723, 2724, 2725, 2726, 2727, 2728, 2729, 2730, 2731, 2732, 2733, 2734, 2735, 2736, 2737, 2738, 2739, 2740, 2741, 2742, 2743, 2744, 2745, 2746, 2747, 2748, 2749, 2750, 2751, 2752, 2753, 2754, 2755, 2756, 2757, 2758, 2759, 2760, 2761, 2762, 2763, 2764, 2765, 2766, 2767, 2768, 2769, 2770, 2771, 2772, 2773, 2774, 2775, 2776, 2777, 2778, 2779, 2780, 2781, 2782, 2783, 2784, 2785, 2786, 2787, 2788, 2789, 2790, 2791, 2792, 2793, 2794, 2795, 2796, 2797, 2798, 2799, 2800, 2801, 2802, 2803, 2804, 2805, 2806, 2807, 2808, 2809, 2810, 2811, 2812, 2813, 2814, 2815, 2816, 2817, 2818, 2819, 3592, 3593, 3594, 3595, 3596, 3597, 3598, 3599, 3600, 3601, 3602, 3603, 3604, 3605, 3606, 3607, 3608, 3609, 3610, 3611, 3612, 3613, 3614, 3615, 3616, 3617, 3618, 3619, 3620, 3621, 3622, 3623, 3624, 3625, 3626, 3627, 3628, 3629, 3630, 3631, 3632, 3633, 3634, 3635, 3636, 3637, 3638, 3639, 3640, 3641, 3642, 3643, 3644, 3645, 3646, 3647, 3648, 3649, 3650, 3651, 3652, 3653, 3654, 3655, 3656, 3657, 3658, 3659, 3660, 3661, 3662, 3663, 3664, 3665, 3666, 3667, 3668, 3669, 3670, 3671, 3672, 3673, 3674, 3675, 3676, 3677, 3678, 3679, 3680, 3681, 3682, 3683, 3684, 3685, 3686, 3687, 3688, 3689, 3690, 3691, 3692, 3693, 3694, 3695, 3696, 3697, 3698, 3699, 3700, 3701, 3702, 3703, 3704, 3705, 3706, 3707, 3708, 3709, 3710, 3711, 3712, 3713, 3714, 3715, 3716, 3717, 3718, 3719, 3720, 3721, 3722, 3723, 3724, 3725, 3726, 3727, 3728, 3729, 3730, 3731, 3732, 3733, 3734, 3735, 3736, 3737, 3738, 3739, 3740, 3741, 3742, 3743, 3744, 3745, 3746, 3747, 3748, 3749, 3750, 3751, 3752, 3753, 3754, 3755, 3756, 3757, 3758, 3759, 3760, 3761, 3762, 3763, 3764, 3765, 3766, 3767, 3768, 3769, 3770, 3771, 3772, 3773, 3774, 3775, 3776, 3777, 3778, 3779, 3780, 3781, 3782, 3783, 3784, 3785, 3786, 3787, 3788, 3789, 3790, 3791, 3792, 3793, 3794, 3795, 3796, 3797, 3798, 3799, 3800, 3801, 3802, 3803, 3804, 3805, 3806, 3807, 3808, 3809, 3810, 3811, 3812, 3813, 3814, 3815, 3816, 3817, 3818, 3819, 3820, 3821, 3822, 3823, 3824, 3825, 3826, 3827, 3828, 3829, 3830, 3831, 3832, 3833, 3834, 3835, 3836, 3837, 3838, 3839, 3840, 3841, 3842, 3843, 3844, 3845, 3846, 3847, 4620, 4621, 4622, 4623, 4624, 4625, 4626, 4627, 4628, 4629, 4630, 4631, 4632, 4633, 4634, 4635, 4636, 4637, 4638, 4639, 4640, 4641, 4642, 4643, 4644, 4645, 4646, 4647, 4648, 4649, 4650, 4651, 4652, 4653, 4654, 4655, 4656, 4657, 4658, 4659, 4660, 4661, 4662, 4663, 4664, 4665, 4666, 4667, 4668, 4669, 4670, 4671, 4672, 4673, 4674, 4675, 4676, 4677, 4678, 4679, 4680, 4681, 4682, 4683, 4684, 4685, 4686, 4687, 4688, 4689, 4690, 4691, 4692, 4693, 4694, 4695, 4696, 4697, 4698, 4699, 4700, 4701, 4702, 4703, 4704, 4705, 4706, 4707, 4708, 4709, 4710, 4711, 4712, 4713, 4714, 4715, 4716, 4717, 4718, 4719, 4720, 4721, 4722, 4723, 4724, 4725, 4726, 4727, 4728, 4729, 4730, 4731, 4732, 4733, 4734, 4735, 4736, 4737, 4738, 4739, 4740, 4741, 4742, 4743, 4744, 4745, 4746, 4747, 4748, 4749, 4750, 4751, 4752, 4753, 4754, 4755, 4756, 4757, 4758, 4759, 4760, 4761, 4762, 4763, 4764, 4765, 4766, 4767, 4768, 4769, 4770, 4771, 4772, 4773, 4774, 4775, 4776, 4777, 4778, 4779, 4780, 4781, 4782, 4783, 4784, 4785, 4786, 4787, 4788, 4789, 4790, 4791, 4792, 4793, 4794, 4795, 4796, 4797, 4798, 4799, 4800, 4801, 4802, 4803, 4804, 4805, 4806, 4807, 4808, 4809, 4810, 4811, 4812, 4813, 4814, 4815, 4816, 4817, 4818, 4819, 4820, 4821, 4822, 4823, 4824, 4825, 4826, 4827, 4828, 4829, 4830, 4831, 4832, 4833, 4834, 4835, 4836, 4837, 4838, 4839, 4840, 4841, 4842, 4843, 4844, 4845, 4846, 4847, 4848, 4849, 4850, 4851, 4852, 4853, 4854, 4855, 4856, 4857, 4858, 4859, 4860, 4861, 4862, 4863, 4864, 4865, 4866, 4867, 4868, 4869, 4870, 4871, 4872, 4873, 4874, 4875, 5392, 5393, 5394, 5395, 5396, 5397, 5398, 5399, 5400, 5401, 5402, 5403, 5404, 5405, 5406, 5407, 5408, 5409, 5410, 5411, 5412, 5413, 5414, 5415, 5416, 5417, 5418, 5419, 5420, 5421, 5422, 5423, 5424, 5425, 5426, 5427, 5428, 5429, 5430, 5431, 5432, 5433, 5434, 5435, 5436, 5437, 5438, 5439, 5440, 5441, 5442, 5443, 5444, 5445, 5446, 5447, 5448, 5449, 5450, 5451, 5452, 5453, 5454, 5455, 5456, 5457, 5458, 5459, 5460, 5461, 5462, 5463, 5464, 5465, 5466, 5467, 5468, 5469, 5470, 5471, 5472, 5473, 5474, 5475, 5476, 5477, 5478, 5479, 5480, 5481, 5482, 5483, 5484, 5485, 5486, 5487, 5488, 5489, 5490, 5491, 5492, 5493, 5494, 5495, 5496, 5497, 5498, 5499, 5500, 5501, 5502, 5503, 5504, 5505, 5506, 5507, 5508, 5509, 5510, 5511, 5512, 5513, 5514, 5515, 5516, 5517, 5518, 5519, 5520, 5521, 5522, 5523, 5524, 5525, 5526, 5527, 5528, 5529, 5530, 5531, 5532, 5533, 5534, 5535, 5536, 5537, 5538, 5539, 5540, 5541, 5542, 5543, 5544, 5545, 5546, 5547, 5548, 5549, 5550, 5551, 5552, 5553, 5554, 5555, 5556, 5557, 5558, 5559, 5560, 5561, 5562, 5563, 5564, 5565, 5566, 5567, 5568, 5569, 5570, 5571, 5572, 5573, 5574, 5575, 5576, 5577, 5578, 5579, 5580, 5581, 5582, 5583, 5584, 5585, 5586, 5587, 5588, 5589, 5590, 5591, 5592, 5593, 5594, 5595, 5596, 5597, 5598, 5599, 5600, 5601, 5602, 5603, 5604, 5605, 5606, 5607, 5608, 5609, 5610, 5611, 5612, 5613, 5614, 5615, 5616, 5617, 5618, 5619, 5620, 5621, 5622, 5623, 5624, 5625, 5626, 5627, 5628, 5629, 5630, 5631, 5632, 5633, 5634, 5635, 5636, 5637, 5638, 5639, 5640, 5641, 5642, 5643, 5644, 5645, 5646, 5647, 5908, 5909, 5910, 5911, 5912, 5913, 5914, 5915, 5916, 5917, 5918, 5919, 5920, 5921, 5922, 5923, 5924, 5925, 5926, 5927, 5928, 5929, 5930, 5931, 5932, 5933, 5934, 5935, 5936, 5937, 5938, 5939, 5940, 5941, 5942, 5943, 5944, 5945, 5946, 5947, 5948, 5949, 5950, 5951, 5952, 5953, 5954, 5955, 5956, 5957, 5958, 5959, 5960, 5961, 5962, 5963, 5964, 5965, 5966, 5967, 5968, 5969, 5970, 5971, 5972, 5973, 5974, 5975, 5976, 5977, 5978, 5979, 5980, 5981, 5982, 5983, 5984, 5985, 5986, 5987, 5988, 5989, 5990, 5991, 5992, 5993, 5994, 5995, 5996, 5997, 5998, 5999, 6000, 6001, 6002, 6003, 6004, 6005, 6006, 6007, 6008, 6009, 6010, 6011, 6012, 6013, 6014, 6015, 6016, 6017, 6018, 6019, 6020, 6021, 6022, 6023, 6024, 6025, 6026, 6027, 6028, 6029, 6030, 6031, 6032, 6033, 6034, 6035, 6036, 6037, 6038, 6039, 6040, 6041, 6042, 6043, 6044, 6045, 6046, 6047, 6048, 6049, 6050, 6051, 6052, 6053, 6054, 6055, 6056, 6057, 6058, 6059, 6060, 6061, 6062, 6063, 6064, 6065, 6066, 6067, 6068, 6069, 6070, 6071, 6072, 6073, 6074, 6075, 6076, 6077, 6078, 6079, 6080, 6081, 6082, 6083, 6084, 6085, 6086, 6087, 6088, 6089, 6090, 6091, 6092, 6093, 6094, 6095, 6096, 6097, 6098, 6099, 6100, 6101, 6102, 6103, 6104, 6105, 6106, 6107, 6108, 6109, 6110, 6111, 6112, 6113, 6114, 6115, 6116, 6117, 6118, 6119, 6120, 6121, 6122, 6123, 6124, 6125, 6126, 6127, 6128, 6129, 6130, 6131, 6132, 6133, 6134, 6135, 6136, 6137, 6138, 6139, 6140, 6141, 6142, 6143, 6144, 6145, 6146, 6147, 6148, 6149, 6150, 6151, 6152, 6153, 6154, 6155, 6156, 6157, 6158, 6159, 6160, 6161, 6162, 6163, 6168, 6169, 6170, 6171, 6172, 6173, 6174, 6175, 6176, 6177, 6178, 6179, 6180, 6181, 6182, 6183, 6184, 6185, 6186, 6187, 6188, 6189, 6190, 6191, 6192, 6193, 6194, 6195, 6196, 6197, 6198, 6199, 6200, 6201, 6202, 6203, 6204, 6205, 6206, 6207, 6208, 6209, 6210, 6211, 6212, 6213, 6214, 6215, 6216, 6217, 6218, 6219, 6220, 6221, 6222, 6223, 6224, 6225, 6226, 6227, 6228, 6229, 6230, 6231, 6232, 6233, 6234, 6235, 6236, 6237, 6238, 6239, 6240, 6241, 6242, 6243, 6244, 6245, 6246, 6247, 6248, 6249, 6250, 6251, 6252, 6253, 6254, 6255, 6256, 6257, 6258, 6259, 6260, 6261, 6262, 6263, 6264, 6265, 6266, 6267, 6268, 6269, 6270, 6271, 6272, 6273, 6274, 6275, 6276, 6277, 6278, 6279, 6280, 6281, 6282, 6283, 6284, 6285, 6286, 6287, 6288, 6289, 6290, 6291, 6292, 6293, 6294, 6295, 6296, 6297, 6298, 6299, 6300, 6301, 6302, 6303, 6304, 6305, 6306, 6307, 6308, 6309, 6310, 6311, 6312, 6313, 6314, 6315, 6316, 6317, 6318, 6319, 6320, 6321, 6322, 6323, 6324, 6325, 6326, 6327, 6328, 6329, 6330, 6331, 6332, 6333, 6334, 6335, 6336, 6337, 6338, 6339, 6340, 6341, 6342, 6343, 6344, 6345, 6346, 6347, 6348, 6349, 6350, 6351, 6352, 6353, 6354, 6355, 6356, 6357, 6358, 6359, 6360, 6361, 6362, 6363, 6364, 6365, 6366, 6367, 6368, 6369, 6370, 6371, 6372, 6373, 6374, 6375, 6376, 6377, 6378, 6379, 6380, 6381, 6382, 6383, 6384, 6385, 6386, 6387, 6388, 6389, 6390, 6391, 6392, 6393, 6394, 6395, 6396, 6397, 6398, 6399, 6400, 6401, 6402, 6403, 6404, 6405, 6406, 6407, 6408, 6409, 6410, 6411, 6412, 6413, 6414, 6415, 6416, 6417, 6418, 6419, 6420, 6421, 6422, 6423);
begin

	comp: EntityName generic map (word_size => 8, entries =>6400)
									port map(clk => clk_i, rst => rst_i, en => en_i, go => go_i, done => done_i, readnotwrite => readnotwrite_i, 
									address => address_i, data_in => data_in_i, data_out => data_out_i);

	clk_i <= not(clk_i) after 0.5 ns;
	
	rst_proc : process 
		begin			
			rst_i <= '1';
			wait for 1536 ns;
			rst_i <= '0';
			wait;
	end process;

	cnt_proc: process(rst_i, clk_i) 
		variable cnt : integer := 0;
		variable writeOutputs : integer := 0;
		begin
			if(rst_i = '1') then
				cnt := 0;
			elsif (clk_i'event and clk_i = '1') then
				if (cnt = 6399 and done_i = '0') then
					cnt := 0;
				elsif done_i = '1' then
					cnt := 0;
					writeOutputs := 1;
				else 
					if(writeOutputs /= 1) then
						cnt := cnt + 1;
					else
						cnt := result_address_vector(cnt);
					end if;
				end if;
			end if;
			
			address_i <= std_logic_vector(to_unsigned(cnt, 8));
	end process;

	wrt_proc: process
		variable first : boolean := true;
		begin
			if first then
				wait until en_i'event and en_i = '1' and readnotwrite_i = '0';
				first := false;
			else
				wait until en_i = '1' and readnotwrite_i = '0';
			end if;
			data_in_i <= std_logic_vector(to_unsigned(0, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(2, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(3, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(4, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(5, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(6, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(7, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(8, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(9, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(10, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(11, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(12, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(13, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(14, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(15, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(16, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(17, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(18, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(19, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(20, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(21, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(22, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(23, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(24, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(25, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(26, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(27, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(28, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(29, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(30, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(31, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(32, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(33, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(34, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(35, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(36, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(37, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(38, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(39, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(40, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(41, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(42, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(43, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(44, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(45, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(46, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(47, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(48, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(49, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(50, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(51, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(52, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(53, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(54, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(55, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(56, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(57, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(58, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(59, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(60, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(61, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(62, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(63, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(64, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(65, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(66, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(67, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(68, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(69, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(70, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(71, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(72, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(73, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(74, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(75, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(76, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(77, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(78, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(79, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(80, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(81, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(82, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(83, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(84, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(85, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(86, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(87, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(88, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(89, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(90, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(91, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(92, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(93, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(94, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(95, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(96, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(97, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(98, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(99, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(100, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(101, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(102, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(103, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(104, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(105, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(106, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(107, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(108, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(109, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(110, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(111, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(112, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(113, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(114, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(115, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(116, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(117, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(118, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(119, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(120, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(121, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(122, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(123, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(124, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(125, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(126, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(127, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(128, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(129, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(130, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(131, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(132, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(133, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(134, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(135, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(136, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(137, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(138, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(139, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(140, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(141, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(142, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(143, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(144, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(145, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(146, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(147, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(148, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(149, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(150, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(151, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(152, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(153, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(154, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(155, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(156, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(157, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(158, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(159, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(160, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(161, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(162, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(163, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(164, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(165, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(166, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(167, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(168, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(169, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(170, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(171, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(172, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(173, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(174, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(175, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(176, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(177, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(178, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(179, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(180, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(181, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(182, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(183, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(184, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(185, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(186, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(187, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(188, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(189, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(190, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(191, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(192, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(193, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(194, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(195, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(196, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(197, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(198, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(199, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(200, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(201, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(202, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(203, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(204, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(205, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(206, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(207, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(208, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(209, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(210, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(211, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(212, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(213, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(214, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(215, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(216, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(217, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(218, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(219, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(220, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(221, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(222, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(223, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(224, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(225, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(226, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(227, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(228, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(229, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(230, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(231, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(232, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(233, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(234, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(235, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(236, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(237, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(238, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(239, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(240, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(241, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(242, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(243, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(244, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(245, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(246, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(247, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(248, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(249, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(250, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(251, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(252, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(253, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(254, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(255, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(256, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(257, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(258, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(259, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(260, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(261, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(262, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(263, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(264, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(265, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(266, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(267, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(268, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(269, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(270, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(271, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(272, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(273, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(274, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(275, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(276, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(277, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(278, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(279, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(280, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(281, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(282, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(283, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(284, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(285, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(286, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(287, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(288, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(289, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(290, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(291, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(292, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(293, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(294, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(295, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(296, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(297, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(298, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(299, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(300, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(301, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(302, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(303, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(304, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(305, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(306, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(307, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(308, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(309, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(310, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(311, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(312, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(313, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(314, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(315, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(316, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(317, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(318, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(319, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(320, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(321, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(322, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(323, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(324, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(325, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(326, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(327, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(328, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(329, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(330, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(331, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(332, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(333, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(334, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(335, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(336, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(337, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(338, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(339, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(340, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(341, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(342, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(343, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(344, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(345, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(346, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(347, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(348, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(349, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(350, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(351, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(352, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(353, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(354, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(355, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(356, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(357, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(358, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(359, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(360, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(361, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(362, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(363, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(364, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(365, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(366, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(367, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(368, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(369, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(370, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(371, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(372, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(373, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(374, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(375, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(376, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(377, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(378, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(379, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(380, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(381, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(382, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(383, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(384, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(385, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(386, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(387, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(388, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(389, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(390, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(391, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(392, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(393, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(394, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(395, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(396, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(397, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(398, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(399, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(400, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(401, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(402, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(403, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(404, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(405, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(406, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(407, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(408, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(409, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(410, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(411, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(412, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(413, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(414, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(415, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(416, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(417, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(418, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(419, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(420, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(421, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(422, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(423, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(424, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(425, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(426, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(427, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(428, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(429, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(430, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(431, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(432, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(433, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(434, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(435, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(436, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(437, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(438, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(439, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(440, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(441, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(442, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(443, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(444, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(445, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(446, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(447, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(448, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(449, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(450, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(451, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(452, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(453, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(454, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(455, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(456, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(457, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(458, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(459, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(460, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(461, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(462, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(463, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(464, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(465, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(466, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(467, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(468, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(469, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(470, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(471, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(472, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(473, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(474, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(475, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(476, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(477, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(478, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(479, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(480, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(481, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(482, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(483, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(484, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(485, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(486, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(487, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(488, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(489, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(490, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(491, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(492, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(493, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(494, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(495, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(496, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(497, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(498, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(499, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(500, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(501, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(502, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(503, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(504, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(505, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(506, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(507, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(508, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(509, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(510, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(511, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(512, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(513, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(514, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(515, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(516, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(517, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(518, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(519, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(520, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(521, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(522, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(523, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(524, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(525, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(526, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(527, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(528, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(529, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(530, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(531, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(532, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(533, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(534, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(535, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(536, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(537, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(538, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(539, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(540, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(541, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(542, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(543, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(544, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(545, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(546, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(547, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(548, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(549, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(550, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(551, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(552, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(553, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(554, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(555, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(556, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(557, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(558, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(559, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(560, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(561, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(562, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(563, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(564, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(565, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(566, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(567, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(568, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(569, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(570, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(571, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(572, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(573, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(574, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(575, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(576, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(577, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(578, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(579, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(580, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(581, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(582, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(583, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(584, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(585, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(586, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(587, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(588, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(589, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(590, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(591, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(592, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(593, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(594, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(595, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(596, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(597, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(598, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(599, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(600, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(601, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(602, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(603, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(604, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(605, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(606, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(607, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(608, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(609, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(610, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(611, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(612, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(613, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(614, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(615, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(616, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(617, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(618, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(619, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(620, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(621, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(622, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(623, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(624, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(625, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(626, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(627, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(628, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(629, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(630, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(631, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(632, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(633, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(634, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(635, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(636, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(637, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(638, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(639, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(640, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(641, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(642, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(643, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(644, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(645, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(646, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(647, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(648, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(649, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(650, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(651, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(652, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(653, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(654, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(655, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(656, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(657, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(658, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(659, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(660, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(661, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(662, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(663, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(664, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(665, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(666, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(667, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(668, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(669, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(670, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(671, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(672, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(673, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(674, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(675, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(676, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(677, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(678, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(679, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(680, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(681, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(682, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(683, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(684, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(685, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(686, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(687, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(688, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(689, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(690, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(691, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(692, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(693, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(694, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(695, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(696, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(697, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(698, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(699, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(700, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(701, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(702, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(703, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(704, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(705, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(706, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(707, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(708, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(709, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(710, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(711, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(712, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(713, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(714, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(715, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(716, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(717, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(718, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(719, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(720, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(721, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(722, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(723, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(724, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(725, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(726, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(727, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(728, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(729, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(730, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(731, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(732, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(733, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(734, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(735, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(736, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(737, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(738, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(739, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(740, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(741, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(742, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(743, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(744, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(745, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(746, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(747, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(748, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(749, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(750, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(751, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(752, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(753, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(754, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(755, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(756, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(757, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(758, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(759, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(760, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(761, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(762, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(763, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(764, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(765, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(766, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(767, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(768, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(769, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(770, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(771, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(772, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(773, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(774, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(775, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(776, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(777, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(778, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(779, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(780, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(781, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(782, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(783, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(784, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(785, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(786, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(787, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(788, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(789, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(790, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(791, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(792, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(793, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(794, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(795, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(796, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(797, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(798, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(799, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(800, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(801, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(802, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(803, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(804, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(805, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(806, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(807, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(808, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(809, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(810, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(811, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(812, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(813, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(814, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(815, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(816, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(817, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(818, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(819, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(820, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(821, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(822, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(823, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(824, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(825, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(826, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(827, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(828, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(829, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(830, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(831, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(832, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(833, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(834, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(835, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(836, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(837, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(838, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(839, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(840, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(841, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(842, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(843, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(844, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(845, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(846, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(847, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(848, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(849, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(850, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(851, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(852, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(853, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(854, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(855, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(856, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(857, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(858, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(859, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(860, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(861, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(862, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(863, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(864, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(865, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(866, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(867, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(868, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(869, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(870, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(871, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(872, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(873, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(874, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(875, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(876, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(877, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(878, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(879, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(880, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(881, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(882, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(883, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(884, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(885, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(886, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(887, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(888, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(889, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(890, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(891, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(892, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(893, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(894, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(895, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(896, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(897, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(898, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(899, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(900, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(901, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(902, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(903, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(904, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(905, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(906, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(907, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(908, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(909, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(910, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(911, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(912, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(913, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(914, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(915, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(916, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(917, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(918, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(919, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(920, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(921, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(922, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(923, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(924, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(925, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(926, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(927, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(928, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(929, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(930, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(931, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(932, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(933, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(934, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(935, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(936, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(937, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(938, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(939, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(940, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(941, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(942, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(943, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(944, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(945, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(946, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(947, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(948, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(949, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(950, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(951, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(952, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(953, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(954, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(955, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(956, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(957, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(958, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(959, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(960, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(961, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(962, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(963, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(964, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(965, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(966, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(967, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(968, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(969, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(970, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(971, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(972, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(973, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(974, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(975, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(976, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(977, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(978, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(979, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(980, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(981, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(982, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(983, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(984, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(985, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(986, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(987, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(988, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(989, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(990, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(991, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(992, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(993, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(994, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(995, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(996, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(997, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(998, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(999, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1000, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1001, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1002, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1003, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1004, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1005, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1006, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1007, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1008, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1009, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1010, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1011, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1012, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1013, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1014, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1015, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1016, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1017, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1018, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1019, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1020, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1021, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1022, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1023, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1024, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1025, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1026, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1027, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1028, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1029, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1030, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1031, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1032, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1033, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1034, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1035, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1036, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1037, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1038, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1039, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1040, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1041, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1042, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1043, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1044, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1045, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1046, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1047, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1048, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1049, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1050, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1051, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1052, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1053, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1054, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1055, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1056, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1057, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1058, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1059, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1060, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1061, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1062, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1063, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1064, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1065, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1066, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1067, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1068, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1069, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1070, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1071, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1072, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1073, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1074, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1075, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1076, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1077, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1078, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1079, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1080, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1081, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1082, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1083, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1084, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1085, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1086, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1087, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1088, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1089, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1090, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1091, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1092, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1093, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1094, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1095, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1096, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1097, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1098, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1099, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1100, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1101, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1102, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1103, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1104, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1105, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1106, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1107, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1108, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1109, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1110, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1111, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1112, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1113, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1114, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1115, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1116, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1117, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1118, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1119, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1120, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1121, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1122, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1123, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1124, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1125, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1126, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1127, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1128, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1129, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1130, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1131, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1132, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1133, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1134, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1135, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1136, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1137, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1138, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1139, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1140, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1141, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1142, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1143, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1144, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1145, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1146, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1147, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1148, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1149, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1150, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1151, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1152, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1153, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1154, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1155, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1156, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1157, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1158, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1159, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1160, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1161, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1162, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1163, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1164, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1165, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1166, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1167, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1168, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1169, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1170, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1171, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1172, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1173, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1174, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1175, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1176, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1177, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1178, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1179, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1180, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1181, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1182, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1183, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1184, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1185, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1186, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1187, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1188, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1189, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1190, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1191, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1192, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1193, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1194, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1195, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1196, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1197, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1198, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1199, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1200, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1201, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1202, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1203, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1204, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1205, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1206, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1207, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1208, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1209, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1210, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1211, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1212, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1213, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1214, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1215, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1216, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1217, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1218, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1219, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1220, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1221, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1222, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1223, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1224, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1225, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1226, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1227, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1228, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1229, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1230, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1231, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1232, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1233, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1234, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1235, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1236, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1237, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1238, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1239, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1240, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1241, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1242, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1243, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1244, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1245, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1246, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1247, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1248, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1249, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1250, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1251, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1252, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1253, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1254, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1255, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1256, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1257, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1258, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1259, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1260, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1261, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1262, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1263, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1264, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1265, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1266, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1267, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1268, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1269, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1270, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1271, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1272, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1273, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1274, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1275, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1276, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1277, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1278, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1279, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1280, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1281, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1282, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1283, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1284, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1285, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1286, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1287, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1288, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1289, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1290, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1291, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1292, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1293, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1294, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1295, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1296, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1297, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1298, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1299, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1300, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1301, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1302, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1303, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1304, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1305, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1306, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1307, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1308, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1309, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1310, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1311, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1312, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1313, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1314, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1315, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1316, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1317, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1318, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1319, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1320, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1321, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1322, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1323, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1324, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1325, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1326, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1327, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1328, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1329, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1330, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1331, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1332, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1333, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1334, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1335, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1336, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1337, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1338, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1339, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1340, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1341, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1342, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1343, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1344, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1345, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1346, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1347, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1348, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1349, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1350, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1351, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1352, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1353, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1354, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1355, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1356, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1357, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1358, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1359, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1360, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1361, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1362, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1363, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1364, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1365, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1366, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1367, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1368, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1369, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1370, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1371, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1372, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1373, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1374, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1375, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1376, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1377, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1378, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1379, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1380, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1381, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1382, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1383, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1384, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1385, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1386, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1387, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1388, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1389, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1390, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1391, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1392, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1393, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1394, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1395, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1396, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1397, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1398, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1399, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1400, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1401, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1402, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1403, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1404, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1405, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1406, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1407, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1408, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1409, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1410, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1411, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1412, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1413, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1414, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1415, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1416, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1417, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1418, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1419, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1420, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1421, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1422, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1423, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1424, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1425, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1426, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1427, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1428, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1429, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1430, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1431, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1432, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1433, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1434, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1435, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1436, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1437, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1438, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1439, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1440, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1441, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1442, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1443, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1444, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1445, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1446, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1447, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1448, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1449, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1450, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1451, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1452, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1453, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1454, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1455, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1456, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1457, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1458, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1459, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1460, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1461, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1462, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1463, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1464, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1465, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1466, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1467, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1468, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1469, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1470, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1471, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1472, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1473, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1474, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1475, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1476, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1477, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1478, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1479, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1480, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1481, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1482, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1483, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1484, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1485, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1486, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1487, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1488, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1489, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1490, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1491, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1492, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1493, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1494, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1495, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1496, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1497, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1498, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1499, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1500, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1501, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1502, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1503, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1504, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1505, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1506, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1507, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1508, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1509, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1510, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1511, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1512, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1513, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1514, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1515, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1516, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1517, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1518, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1519, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1520, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1521, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1522, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1523, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1524, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1525, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1526, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1527, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1528, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1529, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1530, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1531, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1532, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1533, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1534, 8));
			wait for 1 ns;		
			data_in_i <= std_logic_vector(to_unsigned(1535, 8));
			wait for 1 ns;		
	end process;

	en_proc: process	
		variable first : boolean := true;
		begin
			if first then
				wait for 1536 ns;
				first := false;
			end if;
			en_i <= '1';
			readnotwrite_i <= '0';
			wait for 1536 ns;
			en_i <= '0';
			wait until done_i'event and done_i = '0';
			en_i <= '1';
			readnotwrite_i <= '1';
			wait for 1536 ns;
	end process;

	go_proc: process
		begin
			wait until en_i'event and en_i = '0';
			go_i <= '1';
			wait for 1 ns;
			go_i <= '0';	
	end process;


end test;